LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Decod7Seg IS
	PORT(e:IN STD_LOGIC_VECTOR(3 downto 0);
		  s:OUT STD_LOGIC_VECTOR(6 downto 0));
END ENTITY;

ARCHITECTURE bhv OF Decod7Seg IS
BEGIN
	WITH e SELECT
	  	 s <= "1000000" WHEN "0000",
				"1111001" WHEN "0001",
				"0100100" WHEN "0010",
				"0110000" WHEN "0011",
				"0011001" WHEN "0100",
				"0010010" WHEN "0101",
				"0000010" WHEN "0110",
				"0111000" WHEN "0111",
				"0000000" WHEN "1000",
				"0010000" WHEN "1001",
				"1111111" WHEN OTHERS;
END ARCHITECTURE;
